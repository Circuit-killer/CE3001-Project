module CPU(Clk, Rst);
  
  input Clk, Rst;
  
  //reg Buff[]
  
endmodule
            
